library verilog;
use verilog.vl_types.all;
entity HALF_ADDSUB_vlg_vec_tst is
end HALF_ADDSUB_vlg_vec_tst;
